`ifndef UARTBASETESTPKG_INCLUDED_
`define UARTBASETESTPKG_INCLUDED_
//--------------------------------------------------------------------------------------------
// Package:UartBaseTestPkg
//--------------------------------------------------------------------------------------------
package UartBaseTestPkg;
  `include "uvm_macros.svh"
  
  //-------------------------------------------------------
  // Import uvm package
  //-------------------------------------------------------
  import uvm_pkg :: *;
  import UartGlobalPkg :: *;

  //-------------------------------------------------------
  // Importing the required packages
  //-------------------------------------------------------
  import UartTxPkg ::*;
  import UartRxPkg :: *;
  import UartEnvPkg :: *;
  import UartTxSequencePkg :: *;
  import UartRxSequencePkg :: *;
  import UartVirtualSequencePkg::*;
  
  //including base_test for testing
  
  `include "UartBaseTest.sv"
  `include "UartEvenParityTest.sv"
  `include "UartOddParityTest.sv"


  `include "UartSample13BaudRate4800Datatype5EvenParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype5EvenParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype5OddParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype5OddParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype6EvenParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype6EvenParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype6OddParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype6OddParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype7EvenParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype7EvenParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype7OddParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype7OddParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype8EvenParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype8EvenParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype8OddParityStopbit1.sv"
  `include "UartSample13BaudRate4800Datatype8OddParityStopbit2.sv"
  `include "UartSample13BaudRate4800Datatype8EvenParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype5EvenParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype5EvenParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype5OddParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype5OddParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype6EvenParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype6EvenParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype6OddParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype6OddParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype7EvenParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype7EvenParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype7OddParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype7OddParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype8EvenParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype8EvenParityStopbit2.sv"
  `include "UartSample13BaudRate9600Datatype8OddParityStopbit1.sv"
  `include "UartSample13BaudRate9600Datatype8OddParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype5EvenParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype5EvenParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype5OddParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype5OddParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype6EvenParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype6EvenParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype6OddParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype6OddParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype7EvenParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype7EvenParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype7OddParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype7OddParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype8EvenParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype8EvenParityStopbit2.sv"
  `include "UartSample13BaudRate19200Datatype8OddParityStopbit1.sv"
  `include "UartSample13BaudRate19200Datatype8OddParityStopbit2.sv"
  `include "UartSample16BaudRate4800Datatype5EvenParityStopbit1.sv"
  `include "UartSample16BaudRate9600Datatype7EvenParityStopbit1.sv"
  `include "UartSample16BaudRate9600Datatype7EvenParityStopbit2.sv"
  `include "UartSample16BaudRate9600Datatype7OddParityStopbit1.sv"
  `include "UartSample16BaudRate9600Datatype7OddParityStopbit2.sv"
  `include "UartSample16BaudRate9600Datatype8EvenParityStopbit1.sv"
  `include "UartSample16BaudRate9600Datatype8EvenParityStopbit2.sv"
  `include "UartSample16BaudRate9600Datatype8OddParityStopbit1.sv"
  `include "UartSample16BaudRate9600Datatype8OddParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype5EvenParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype5EvenParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype5OddParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype5OddParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype6EvenParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype6EvenParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype6OddParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype6OddParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype7EvenParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype7EvenParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype7OddParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype7OddParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype8EvenParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype8EvenParityStopbit2.sv"
  `include "UartSample16BaudRate19200Datatype8OddParityStopbit1.sv"
  `include "UartSample16BaudRate19200Datatype8OddParityStopbit2.sv"

  //  No Parity Test cases

  `include UartSample13BaudRate19200Datatype5NoParityStopbit1.sv
  `include UartSample13BaudRate19200Datatype5NoParityStopbit2.sv
  `include UartSample13BaudRate19200Datatype6NoParityStopbit1.sv
  `include UartSample13BaudRate19200Datatype6NoParityStopbit2.sv
  `include UartSample13BaudRate19200Datatype7NoParityStopbit1.sv
  `include UartSample13BaudRate19200Datatype7NoParityStopbit2.sv
  `include UartSample13BaudRate19200Datatype8NoParityStopbit1.sv
  `include UartSample13BaudRate19200Datatype8NoParityStopbit2.sv
  `include UartSample13BaudRate4800Datatype5NoParityStopbit1.sv
  `include UartSample13BaudRate4800Datatype5NoParityStopbit2.sv
  `include UartSample13BaudRate4800Datatype6NoParityStopbit1.sv
  `include UartSample13BaudRate4800Datatype6NoParityStopbit2.sv
  `include UartSample13BaudRate4800Datatype7NoParityStopbit1.sv
  `include UartSample13BaudRate4800Datatype7NoParityStopbit2.sv
  `include UartSample13BaudRate4800Datatype8NoParityStopbit1.sv
  `include UartSample13BaudRate4800Datatype8NoParityStopbit2.sv
  `include UartSample13BaudRate9600Datatype5NoParityStopbit1.sv
  `include UartSample13BaudRate9600Datatype5NoParityStopbit2.sv
  `include UartSample13BaudRate9600Datatype6NoParityStopbit1.sv
  `include UartSample13BaudRate9600Datatype6NoParityStopbit2.sv
  `include UartSample13BaudRate9600Datatype7NoParityStopbit1.sv
  `include UartSample13BaudRate9600Datatype7NoParityStopbit2.sv
  `include UartSample13BaudRate9600Datatype8NoParityStopbit1.sv
  `include UartSample13BaudRate9600Datatype8NoParityStopbit2.sv
  `include UartSample16BaudRate19200Datatype5NoParityStopbit1.sv
  `include UartSample16BaudRate19200Datatype5NoParityStopbit2.sv
  `include UartSample16BaudRate19200Datatype6NoParityStopbit1.sv
  `include UartSample16BaudRate19200Datatype6NoParityStopbit2.sv
  `include UartSample16BaudRate19200Datatype7NoParityStopbit1.sv
  `include UartSample16BaudRate19200Datatype7NoParityStopbit2.sv
  `include UartSample16BaudRate19200Datatype8NoParityStopbit1.sv
  `include UartSample16BaudRate19200Datatype8NoParityStopbit2.sv
  `include UartSample16BaudRate4800Datatype5NoParityStopbit1.sv
  `include UartSample16BaudRate4800Datatype5NoParityStopbit2.sv
  `include UartSample16BaudRate4800Datatype6NoParityStopbit1.sv
  `include UartSample16BaudRate4800Datatype6NoParityStopbit2.sv
  `include UartSample16BaudRate4800Datatype7NoParityStopbit1.sv
  `include UartSample16BaudRate4800Datatype7NoParityStopbit2.sv
  `include UartSample16BaudRate4800Datatype8NoParityStopbit1.sv
  `include UartSample16BaudRate4800Datatype8NoParityStopbit2.sv
  `include UartSample16BaudRate9600Datatype5NoParityStopbit1.sv
  `include UartSample16BaudRate9600Datatype5NoParityStopbit2.sv
  `include UartSample16BaudRate9600Datatype6NoParityStopbit1.sv
  `include UartSample16BaudRate9600Datatype6NoParityStopbit2.sv
  `include UartSample16BaudRate9600Datatype7NoParityStopbit1.sv
  `include UartSample16BaudRate9600Datatype7NoParityStopbit2.sv
  `include UartSample16BaudRate9600Datatype8NoParityStopbit1.sv
  `include UartSample16BaudRate9600Datatype8NoParityStopbit2.sv
  
  //   Error Test cases  
  `include "UartBreakingErrorTest.sv"
  `include "UartEvenParityWithErrorTest.sv"
  `include "UartOddParityWithErrorTest.sv"
  `include "UartFramingErrorEvenParityTest.sv"
endpackage : UartBaseTestPkg
`endif
