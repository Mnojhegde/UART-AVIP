//-------------------------------------------------------
// Importing Uart global package
//-------------------------------------------------------
import UartGlobalPkg::*;

//--------------------------------------------------------------------------------------------
// Interface : UartTxMonitorBfm
//  Connects the master monitor bfm with the master monitor prox
//--------------------------------------------------------------------------------------------

interface UartTxMonitorBfm (input  bit   clk,
                            input  bit   reset,
                            input  bit   tx
                           );

  //-------------------------------------------------------
  // Importing uvm package file
  //-------------------------------------------------------
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  //-------------------------------------------------------
  // Importing the Transmitter package file
  //-------------------------------------------------------
  //import UartTxPkg:: UartTxMonitorProxy;
  
  //Variable: name
  //Used to store the name of the interface

  string name = "UART_TRANSMITTER_MONITOR_BFM"; 

  //Variable: bclk
  //baud clock for uart transmisson/reception
	
  bit bclk;
   
   //Variable: baudRate
  //Used to sample the uart data
	
 // reg[31:0] baudRate = 9600;
  
   //Variable: baudRate
  // Counter to keep track of clock cycles
	
  reg [15:0] counter;  
  
   //Variable: baudDivider
  //to Calculate baud rate divider
	
  reg [15:0] baudDivider;
	

 //Creating the handle for the proxy_driver

 // UartTxMonitorProxy uartTxMonitorProxy;
   

  //-------------------------------------------------------
  // Used to display the name of the interface
  //-------------------------------------------------------
  initial begin
    `uvm_info(name, $sformatf(name),UVM_LOW)
  end

  
  //------------------------------------------------------------------
  // Task: Baud_div
  // this task will calculate the baud divider based on sys clk frequency
  //-------------------------------------------------------------------
  task Baud_div(input oversamplingmethod,input baudrate);
      real clkPeriodStartTime; 
      real clkPeriodStopTime;
      real clkPeriod;
      real clkFrequency;
      int baudDivisor;
      @(posedge clk);
      clkPeriodStartTime = $realtime;
      @(posedge clk);
      clkPeriodStopTime = $realtime; 
      clkPeriod = clkPeriodStopTime - clkPeriodStartTime;
      clkFrequency = ( 10 **9 )/ clkPeriod;

      baudDivisor = (clkFrequency)/(oversamplingmethod * baudrate); 

      BaudClkGenerator(baudDivisor);
    endtask

  //------------------------------------------------------------------
  // Task: BaudClkGenerator
  // this task will generate baud clk based on baud divider
  //-------------------------------------------------------------------

    task BaudClkGenerator(input int baudDivisor);
      static int count=0;
      forever begin 
        @(posedge clk or negedge clk)
    
        if(count == (baudDivisor-1))begin 
          count <= 0;
          baudClk <= ~baudClk;
        end 
        else begin 
          count <= count +1;
        end   
      end
    endtask
	
  //-------------------------------------------------------
  // Task: WaitForReset
  //  Waiting for the system reset
  //-------------------------------------------------------

  task WaitForReset();
    
  endtask: WaitForReset
  

endinterface : UartTxMonitorBfm
