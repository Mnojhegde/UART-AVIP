import UartGlobalPkg::*;
//--------------------------------------------------------------------------------------------
// Interface : UartTxMonitorBfm
//  Connects the master monitor bfm with the master monitor prox
//--------------------------------------------------------------------------------------------
interface UartTxMonitorBfm (input  logic   clk,
                            input  logic reset,
                            input  logic   tx
                           );
  //-------------------------------------------------------
  // Importing uvm package file
  //-------------------------------------------------------
  import uvm_pkg::*;
  `include "uvm_macros.svh"
	
  string name = "UART_TRANSMITTER_MONITOR_BFM";
	
  //Variable: bclk
  //baud clock for uart transmisson/reception
	bit baudClk;

	logic [DATA_WIDTH+2 : 0]concatData;
	int numOfZeroes;
	int breakZeroCount;

	// enum variable for transfer states
	UartTransmitterStateEnum uartTransmitterState;
	
  //-------------------------------------------------------
  // Used to display the name of the interface
  //-------------------------------------------------------
  initial begin
    `uvm_info(name, $sformatf(name),UVM_LOW)
  end

  //------------------------------------------------------------------
  // Task: Baud_div
  // this task will calculate the baud divider based on sys clk frequency
  //-------------------------------------------------------------------
  task GenerateBaudClk(inout UartConfigStruct uartConfigStruct);
      real clkPeriodStartTime;
      real clkPeriodStopTime;
      real clkPeriod;
      real clkFrequency;
      int baudDivisor;
      @(posedge clk);
      clkPeriodStartTime = $realtime;
      @(posedge clk);
      clkPeriodStopTime = $realtime;
      clkPeriod = clkPeriodStopTime - clkPeriodStartTime;
      clkFrequency = ( 10 **9 )/ clkPeriod;
      if(uartConfigStruct.OverSampledBaudFrequencyClk==1)begin
      baudDivisor = (clkFrequency)/(uartConfigStruct.uartOverSamplingMethod * uartConfigStruct.uartBaudRate);
      end
      else begin
      baudDivisor = (clkFrequency)/(uartConfigStruct.uartBaudRate);
      end
      BaudClkGenerator(baudDivisor);
    endtask
	
  //------------------------------------------------------------------
  // Task: BaudClkGenerator
  // this task will generate baud clk based on baud divider
  //-------------------------------------------------------------------
    task BaudClkGenerator(input int baudDiv);
      static int count=0;
      forever begin
        @(posedge clk or negedge clk)
        if(count == (baudDiv-1))begin
          count <= 0;
          baudClk <= ~baudClk;
        end
        else begin
          count <= count +1;
        end
      end
    endtask
	
  //-------------------------------------------------------
  // Task: WaitForReset
  //  Waiting for the system reset
  //-------------------------------------------------------
  task WaitForReset();
    @(negedge reset);
    `uvm_info(name, $sformatf("system reset activated"), UVM_LOW)
		uartTransmitterState = RESET;
    @(posedge reset);
    `uvm_info(name, $sformatf("system reset deactivated"), UVM_LOW)
	  uartTransmitterState = IDLE;
  endtask: WaitForReset
	
	task StartMonitoring(inout UartTxPacketStruct uartTxPacketStruct , inout UartConfigStruct uartConfigStruct);
		Deserializer(uartTxPacketStruct,uartConfigStruct);
  endtask

	function evenParityCompute(input UartConfigStruct uartConfigStruct,input UartTxPacketStruct uartTxPacketStruct);
	  bit parity;
	  case(uartConfigStruct.uartDataType)
	    FIVE_BIT: parity = ^(uartTxPacketStruct.transmissionData[4:0]);
	    SIX_BIT :parity = ^(uartTxPacketStruct.transmissionData[5:0]);
	    SEVEN_BIT: parity = ^(uartTxPacketStruct.transmissionData[6:0]);
	    EIGHT_BIT : parity = ^(uartTxPacketStruct.transmissionData[7:0]);
	  endcase
	return parity;
	endfunction
	function oddParityCompute(input UartConfigStruct uartConfigStruct,input UartTxPacketStruct uartTxPacketStruct);
	  bit parity;
	  case(uartConfigStruct.uartDataType)
	      FIVE_BIT: parity = ~^(uartTxPacketStruct.transmissionData[4:0]);
	      SIX_BIT :parity = ~^(uartTxPacketStruct.transmissionData[5:0]);
	      SEVEN_BIT: parity = ~^(uartTxPacketStruct.transmissionData[6:0]);
	      EIGHT_BIT : parity = ~^(uartTxPacketStruct.transmissionData[7:0]);
	  endcase
	return parity;
	endfunction
	
  //-------------------------------------------------------
  // Task: DeSerializer
  //  converts serial data to parallel
  //-------------------------------------------------------
  task Deserializer(inout UartTxPacketStruct uartTxPacketStruct, inout UartConfigStruct uartConfigStruct);
		// sampling start bit 
	  @(negedge tx);
        if(uartConfigStruct.OverSampledBaudFrequencyClk==1)begin
        	repeat(uartConfigStruct.uartOverSamplingMethod/2) @(posedge baudClk); 
					uartTransmitterState = STARTBIT;
					concatData={concatData,tx};
	

					// sampling data bits 
					for( int i=0 ; i < uartConfigStruct.uartDataType ; i++) begin
          	repeat(uartConfigStruct.uartOverSamplingMethod) @(posedge baudClk); begin
						uartTxPacketStruct.transmissionData[i] = tx;
			      concatData={concatData,tx};
						uartTransmitterState = UartTransmitterStateEnum'(i+3);
          end
        end

				// sampling parity bit 
        if(uartConfigStruct.uartParityEnable ==1) begin
        	repeat(uartConfigStruct.uartOverSamplingMethod) @(posedge baudClk);
					$display("PARITY IS ASSSIGNED AT %t",$time);
					uartTxPacketStruct.parity = tx;
					concatData={concatData,tx};
					uartTransmitterState = PARITYBIT;
					parityCheck(uartConfigStruct,uartTxPacketStruct,tx);
      	end
		$display("OUTSIDE PARITY GEN IS %t",$time);
				// sampling stop bit	
        repeat(uartConfigStruct.uartOverSamplingMethod) @(posedge baudClk);
					concatData={concatData,tx};
					stopBitCheck(uartTxPacketStruct,uartConfigStruct,tx);
					$display("STOP BIT IS BEING ASSIGNED IN  MONITOR AT %t",$time);
					numOfZeroes=$countones(~(concatData));
					breakZeroCount=uartConfigStruct.uartParityEnable ? (uartConfigStruct.uartDataType)+3 :(uartConfigStruct.uartDataType)+2;
					$display("THE NUMBER OF ZEROES IS %0d",numOfZeroes);
					if(numOfZeroes == breakZeroCount)
						uartTxPacketStruct.breakingError =1;
				  else 
						uartTxPacketStruct.breakingError =0;


					$display("THE BREAKING ERROR IS %b",uartTxPacketStruct.breakingError);
					concatData = 'b x;
					numOfZeroes =0;
					uartTransmitterState = IDLE;
					repeat(uartConfigStruct.uartOverSamplingMethod/2) @(posedge baudClk);
					
        end
		
        else if(uartConfigStruct.OverSampledBaudFrequencyClk==0)begin
					// sampling start bit 
					repeat(1)@(posedge baudClk);
					uartTransmitterState = STARTBIT;
					
					// sampling data bits 
					for( int i=0 ; i < uartConfigStruct.uartDataType ; i++) begin
          	@(posedge baudClk)begin
		  				uartTxPacketStruct.transmissionData[i] = tx;
							uartTransmitterState = UartTransmitterStateEnum'(i+3);
        		end
        	end

					// sampling parity bit 
					if(uartConfigStruct.uartParityEnable ==1) begin
        		@(posedge baudClk)
         		uartTxPacketStruct.parity = tx;
						uartTransmitterState = PARITYBIT;
		 				parityCheck(uartConfigStruct,uartTxPacketStruct,tx);
        	end

					// sampling stop bit	
        	@(posedge baudClk);
					uartTransmitterState = STOPBIT;
		      stopBitCheck(uartTxPacketStruct,uartConfigStruct,tx);
      	end
    endtask
	
	task stopBitCheck (inout  UartTxPacketStruct uartTxPacketStruct,input UartConfigStruct uartConfigStruct,input bit tx);
			if (tx == 1) begin
				uartTxPacketStruct.framingError = 0;
				uartTransmitterState = STOPBIT;
			end
			else begin
				uartTxPacketStruct.framingError = 1;
				uartTransmitterState = INVALIDSTOPBIT;
				repeat(uartConfigStruct.uartOverSamplingMethod)@(posedge baudClk);
			end
  	endtask
		
		task parityCheck(inout UartConfigStruct uartConfigStruct,inout UartTxPacketStruct uartTxPacketStruct,input bit tx);
   		int cal_parity;
   		if(uartConfigStruct.uartParityType == EVEN_PARITY)begin
      	cal_parity = evenParityCompute(uartConfigStruct,uartTxPacketStruct);
     	end
      else begin
      	cal_parity = oddParityCompute(uartConfigStruct,uartTxPacketStruct);
      end
			if(tx==cal_parity)begin
      	uartTxPacketStruct.parityError=0;
     	end
     	else begin
     		uartTxPacketStruct.parityError=1;
     	end
  	endtask:parityCheck
endinterface : UartTxMonitorBfm
