class master_monitor_proxy extends uvm_component;
  
  
  `uvm_component_utils(master_monitor_proxy)
  
  master_agent_config master_agent_cfg_h;

  //declaring analysis port for the monitor port
  uvm_analysis_port #(master_tx)master_analysis_port;
  
  //-------------------------------------------------------
  // Externally defined Tasks and Functions
  //-------------------------------------------------------
  extern function new(string name = "master_monitor_proxy", uvm_component parent = null);
  extern function void build_phase(uvm_phase phase);
  extern function void connect_phase(uvm_phase phase);
  extern function void end_of_elaboration_phase(uvm_phase phase);
  extern function void start_of_simulation_phase(uvm_phase phase);
  extern task run_phase(uvm_phase phase);

endclass : master_monitor_proxy

//--------------------------------------------------------------------------------------------
// Construct: new
//--------------------------------------------------------------------------------------------
    function master_monitor_proxy::new(string name = "master_monitor_proxy",
                                 uvm_component parent = null);
  super.new(name, parent);
  
  //creating monitor port
      master_analysis_port=new("master_analysis_port",this);
endfunction : new

//--------------------------------------------------------------------------------------------
// phase - uvm phase
//--------------------------------------------------------------------------------------------
function void master_monitor_proxy::build_phase(uvm_phase phase);
  super.build_phase(phase);
  
  if(!uvm_config_db #(master_agent_config)::get(this,"","master_agent_config",master_agent_cfg_h))begin
    `uvm_fatal("FATAL_master_MONITOR_PROXY_CANNOT_GET_master_AGENT_CONFIG","cannot get() master_agent_cfg_h from uvm_config_db");
  end 

endfunction : build_phase

//--------------------------------------------------------------------------------------------
// Function: connect_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void master_monitor_proxy::connect_phase(uvm_phase phase);
  super.connect_phase(phase);
  
endfunction : connect_phase

//--------------------------------------------------------------------------------------------
// Function: end_of_elaboration_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void master_monitor_proxy::end_of_elaboration_phase(uvm_phase phase);
  super.end_of_elaboration_phase(phase);
endfunction  : end_of_elaboration_phase

//--------------------------------------------------------------------------------------------
// Function: start_of_simulation_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
function void master_monitor_proxy::start_of_simulation_phase(uvm_phase phase);
  super.start_of_simulation_phase(phase);
endfunction : start_of_simulation_phase

//--------------------------------------------------------------------------------------------
// Task: run_phase
// <Description_here>
//
// Parameters:
//  phase - uvm phase
//--------------------------------------------------------------------------------------------
task master_monitor_proxy::run_phase(uvm_phase phase);

  phase.raise_objection(this, "master_monitor_proxy");

  super.run_phase(phase);

  // Work here

  phase.drop_objection(this);

endtask : run_phase
