`ifndef UARTTXASSERTIONTB_INCLUDED_
`define UARTTXASSERTIONTB_INCLUDED_

`include "uvm_macros.svh"
import uvm_pkg :: *;
import UartGlobalPkg :: *;

module UartTxAssertionTb;


endmodule 

`endif
